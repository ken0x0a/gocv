module cv

#include "extra.h"

// enum ColorConversionCodes https://docs.opencv.org/3.4/d8/d01/group__imgproc__color__conversions.html
pub const (
	bgr2_bgra           = 0
	rgb2_rgba           = bgr2_bgra
	bgra2_bgr           = 1
	rgba2_rgb           = bgra2_bgr
	bgr2_rgba           = 2
	rgb2_bgra           = bgr2_rgba
	rgba2_bgr           = 3
	bgra2_rgb           = rgba2_bgr
	bgr2_rgb            = 4
	rgb2_bgr            = bgr2_rgb
	bgra2_rgba          = 5
	rgba2_bgra          = bgra2_rgba
	bgr2_gray           = 6
	rgb2_gray           = 7
	gray2_bgr           = 8
	gray2_rgb           = gray2_bgr
	gray2_bgra          = 9
	gray2_rgba          = gray2_bgra
	bgra2_gray          = 10
	rgba2_gray          = 11
	bgr2_bgr565         = 12
	rgb2_bgr565         = 13
	bgr5652_bgr         = 14
	bgr5652_rgb         = 15
	bgra2_bgr565        = 16
	rgba2_bgr565        = 17
	bgr5652_bgra        = 18
	bgr5652_rgba        = 19
	gray2_bgr565        = 20
	bgr5652_gray        = 21
	bgr2_bgr555         = 22
	rgb2_bgr555         = 23
	bgr5552_bgr         = 24
	bgr5552_rgb         = 25
	bgra2_bgr555        = 26
	rgba2_bgr555        = 27
	bgr5552_bgra        = 28
	bgr5552_rgba        = 29
	gray2_bgr555        = 30
	bgr5552_gray        = 31
	bgr2_xyz            = 32
	rgb2_xyz            = 33
	xyz2_bgr            = 34
	xyz2_rgb            = 35
	bgr2_ycr_cb         = 36
	rgb2_ycr_cb         = 37
	ycr_cb2_bgr         = 38
	ycr_cb2_rgb         = 39
	bgr2_hsv            = 40
	rgb2_hsv            = 41
	bgr2_lab            = 44
	rgb2_lab            = 45
	bgr2_luv            = 50
	rgb2_luv            = 51
	bgr2_hls            = 52
	rgb2_hls            = 53
	hsv2_bgr            = 54
	hsv2_rgb            = 55
	lab2_bgr            = 56
	lab2_rgb            = 57
	luv2_bgr            = 58
	luv2_rgb            = 59
	hls2_bgr            = 60
	hls2_rgb            = 61
	bgr2_hsv_full       = 66
	rgb2_hsv_full       = 67
	bgr2_hls_full       = 68
	rgb2_hls_full       = 69
	hsv2_bgr_full       = 70
	hsv2_rgb_full       = 71
	hls2_bgr_full       = 72
	hls2_rgb_full       = 73
	lbgr2_lab           = 74
	lrgb2_lab           = 75
	lbgr2_luv           = 76
	lrgb2_luv           = 77
	lab2_lbgr           = 78
	lab2_lrgb           = 79
	luv2_lbgr           = 80
	luv2_lrgb           = 81
	bgr2_yuv            = 82
	rgb2_yuv            = 83
	yuv2_bgr            = 84
	yuv2_rgb            = 85
	yuv2_rgb_nv12       = 90
	yuv2_bgr_nv12       = 91
	yuv2_rgb_nv21       = 92
	yuv2_bgr_nv21       = 93
	yuv420sp2_rgb       = yuv2_rgb_nv21
	yuv420sp2_bgr       = yuv2_bgr_nv21
	yuv2_rgba_nv12      = 94
	yuv2_bgra_nv12      = 95
	yuv2_rgba_nv21      = 96
	yuv2_bgra_nv21      = 97
	yuv420sp2_rgba      = yuv2_rgba_nv21
	yuv420sp2_bgra      = yuv2_bgra_nv21
	yuv2_rgb_yv12       = 98
	yuv2_bgr_yv12       = 99
	yuv2_rgb_iyuv       = 100
	yuv2_bgr_iyuv       = 101
	yuv2_rgb_i420       = yuv2_rgb_iyuv
	yuv2_bgr_i420       = yuv2_bgr_iyuv
	yuv420p2_rgb        = yuv2_rgb_yv12
	yuv420p2_bgr        = yuv2_bgr_yv12
	yuv2_rgba_yv12      = 102
	yuv2_bgra_yv12      = 103
	yuv2_rgba_iyuv      = 104
	yuv2_bgra_iyuv      = 105
	yuv2_rgba_i420      = yuv2_rgba_iyuv
	yuv2_bgra_i420      = yuv2_bgra_iyuv
	yuv420p2_rgba       = yuv2_rgba_yv12
	yuv420p2_bgra       = yuv2_bgra_yv12
	yuv2_gray_420       = 106
	yuv2_gray_nv21      = yuv2_gray_420
	yuv2_gray_nv12      = yuv2_gray_420
	yuv2_gray_yv12      = yuv2_gray_420
	yuv2_gray_iyuv      = yuv2_gray_420
	yuv2_gray_i420      = yuv2_gray_420
	yuv420sp2_gray      = yuv2_gray_420
	yuv420p2_gray       = yuv2_gray_420
	yuv2_rgb_uyvy       = 107
	yuv2_bgr_uyvy       = 108
	yuv2_rgb_y422       = yuv2_rgb_uyvy
	yuv2_bgr_y422       = yuv2_bgr_uyvy
	yuv2_rgb_uynv       = yuv2_rgb_uyvy
	yuv2_bgr_uynv       = yuv2_bgr_uyvy
	yuv2_rgba_uyvy      = 111
	yuv2_bgra_uyvy      = 112
	yuv2_rgba_y422      = yuv2_rgba_uyvy
	yuv2_bgra_y422      = yuv2_bgra_uyvy
	yuv2_rgba_uynv      = yuv2_rgba_uyvy
	yuv2_bgra_uynv      = yuv2_bgra_uyvy
	yuv2_rgb_yuy2       = 115
	yuv2_bgr_yuy2       = 116
	yuv2_rgb_yvyu       = 117
	yuv2_bgr_yvyu       = 118
	yuv2_rgb_yuyv       = yuv2_rgb_yuy2
	yuv2_bgr_yuyv       = yuv2_bgr_yuy2
	yuv2_rgb_yunv       = yuv2_rgb_yuy2
	yuv2_bgr_yunv       = yuv2_bgr_yuy2
	yuv2_rgba_yuy2      = 119
	yuv2_bgra_yuy2      = 120
	yuv2_rgba_yvyu      = 121
	yuv2_bgra_yvyu      = 122
	yuv2_rgba_yuyv      = yuv2_rgba_yuy2
	yuv2_bgra_yuyv      = yuv2_bgra_yuy2
	yuv2_rgba_yunv      = yuv2_rgba_yuy2
	yuv2_bgra_yunv      = yuv2_bgra_yuy2
	yuv2_gray_uyvy      = 123
	yuv2_gray_yuy2      = 124
	yuv2_gray_y422      = yuv2_gray_uyvy
	yuv2_gray_uynv      = yuv2_gray_uyvy
	yuv2_gray_yvyu      = yuv2_gray_yuy2
	yuv2_gray_yuyv      = yuv2_gray_yuy2
	yuv2_gray_yunv      = yuv2_gray_yuy2
	rgba2m_rgba         = 125
	m_rgba2_rgba        = 126
	rgb2_yuv_i420       = 127
	bgr2_yuv_i420       = 128
	rgb2_yuv_iyuv       = rgb2_yuv_i420
	bgr2_yuv_iyuv       = bgr2_yuv_i420
	rgba2_yuv_i420      = 129
	bgra2_yuv_i420      = 130
	rgba2_yuv_iyuv      = rgba2_yuv_i420
	bgra2_yuv_iyuv      = bgra2_yuv_i420
	rgb2_yuv_yv12       = 131
	bgr2_yuv_yv12       = 132
	rgba2_yuv_yv12      = 133
	bgra2_yuv_yv12      = 134
	bayer_bg2_bgr       = 46
	bayer_gb2_bgr       = 47
	bayer_rg2_bgr       = 48
	bayer_gr2_bgr       = 49
	bayer_rggb2_bgr     = bayer_bg2_bgr
	bayer_grbg2_bgr     = bayer_gb2_bgr
	bayer_bggr2_bgr     = bayer_rg2_bgr
	bayer_gbrg2_bgr     = bayer_gr2_bgr
	bayer_rggb2_rgb     = bayer_bggr2_bgr
	bayer_grbg2_rgb     = bayer_gbrg2_bgr
	bayer_bggr2_rgb     = bayer_rggb2_bgr
	bayer_gbrg2_rgb     = bayer_grbg2_bgr
	bayer_bg2_rgb       = bayer_rg2_bgr
	bayer_gb2_rgb       = bayer_gr2_bgr
	bayer_rg2_rgb       = bayer_bg2_bgr
	bayer_gr2_rgb       = bayer_gb2_bgr
	bayer_bg2_gray      = 86
	bayer_gb2_gray      = 87
	bayer_rg2_gray      = 88
	bayer_gr2_gray      = 89
	bayer_rggb2_gray    = bayer_bg2_gray
	bayer_grbg2_gray    = bayer_gb2_gray
	bayer_bggr2_gray    = bayer_rg2_gray
	bayer_gbrg2_gray    = bayer_gr2_gray
	bayer_bg2_bgr_vng   = 62
	bayer_gb2_bgr_vng   = 63
	bayer_rg2_bgr_vng   = 64
	bayer_gr2_bgr_vng   = 65
	bayer_rggb2_bgr_vng = bayer_bg2_bgr_vng
	bayer_grbg2_bgr_vng = bayer_gb2_bgr_vng
	bayer_bggr2_bgr_vng = bayer_rg2_bgr_vng
	bayer_gbrg2_bgr_vng = bayer_gr2_bgr_vng
	bayer_rggb2_rgb_vng = bayer_bggr2_bgr_vng
	bayer_grbg2_rgb_vng = bayer_gbrg2_bgr_vng
	bayer_bggr2_rgb_vng = bayer_rggb2_bgr_vng
	bayer_gbrg2_rgb_vng = bayer_grbg2_bgr_vng
	bayer_bg2_rgb_vng   = bayer_rg2_bgr_vng
	bayer_gb2_rgb_vng   = bayer_gr2_bgr_vng
	bayer_rg2_rgb_vng   = bayer_bg2_bgr_vng
	bayer_gr2_rgb_vng   = bayer_gb2_bgr_vng
	bayer_bg2_bgr_ea    = 135
	bayer_gb2_bgr_ea    = 136
	bayer_rg2_bgr_ea    = 137
	bayer_gr2_bgr_ea    = 138
	bayer_rggb2_bgr_ea  = bayer_bg2_bgr_ea
	bayer_grbg2_bgr_ea  = bayer_gb2_bgr_ea
	bayer_bggr2_bgr_ea  = bayer_rg2_bgr_ea
	bayer_gbrg2_bgr_ea  = bayer_gr2_bgr_ea
	bayer_rggb2_rgb_ea  = bayer_bggr2_bgr_ea
	bayer_grbg2_rgb_ea  = bayer_gbrg2_bgr_ea
	bayer_bggr2_rgb_ea  = bayer_rggb2_bgr_ea
	bayer_gbrg2_rgb_ea  = bayer_grbg2_bgr_ea
	bayer_bg2_rgb_ea    = bayer_rg2_bgr_ea
	bayer_gb2_rgb_ea    = bayer_gr2_bgr_ea
	bayer_rg2_rgb_ea    = bayer_bg2_bgr_ea
	bayer_gr2_rgb_ea    = bayer_gb2_bgr_ea
	bayer_bg2_bgra      = 139
	bayer_gb2_bgra      = 140
	bayer_rg2_bgra      = 141
	bayer_gr2_bgra      = 142
	bayer_rggb2_bgra    = bayer_bg2_bgra
	bayer_grbg2_bgra    = bayer_gb2_bgra
	bayer_bggr2_bgra    = bayer_rg2_bgra
	bayer_gbrg2_bgra    = bayer_gr2_bgra
	bayer_rggb2_rgba    = bayer_bggr2_bgra
	bayer_grbg2_rgba    = bayer_gbrg2_bgra
	bayer_bggr2_rgba    = bayer_rggb2_bgra
	bayer_gbrg2_rgba    = bayer_grbg2_bgra
	bayer_bg2_rgba      = bayer_rg2_bgra
	bayer_gb2_rgba      = bayer_gr2_bgra
	bayer_rg2_rgba      = bayer_bg2_bgra
	bayer_gr2_rgba      = bayer_gb2_bgra
	colorcvt_max        = 14
)
