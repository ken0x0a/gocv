module cv
